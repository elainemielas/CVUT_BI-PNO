package CONSCTANS is
	constant COUNTER_WIDTH : integer := 27;
	constant OUTPUT_WIDTH  : integer := 3;
end CONSCTANS;

